///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: tribuf.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::SmartFusion> <Die::A2F200M3F> <Package::484 FBGA>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 
//`timescale <time_units> / <precision>

module tribuf(
input wire a,
input wire en,
output wire b
);
assign b = en? a : 1'bz;
endmodule

