//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Tue Jan 12 13:26:31 2016
// Version: v11.5 SP3 11.5.3.10
//////////////////////////////////////////////////////////////////////

`timescale 1 ns/100 ps

// andor
module andor(
    // Inputs
    SW,
    // Outputs
    LED
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  [1:0] SW;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [5:0] LED;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire         andor_MSS_0_FAB_CLK;
wire   [5:0] LED_0;
wire   [1:0] SW;
wire   [5:0] LED_0_net_0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign LED_0_net_0 = LED_0;
assign LED[5:0]    = LED_0_net_0;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------andor_MSS
andor_MSS andor_MSS_0(
        // Outputs
        .FAB_CLK ( andor_MSS_0_FAB_CLK ) 
        );

//--------myandor
myandor myandor_0(
        // Inputs
        .clk ( andor_MSS_0_FAB_CLK ),
        .SW  ( SW ),
        // Outputs
        .LED ( LED_0 ) 
        );


endmodule
