
module n64_write_command(
    input reg [7:0] command_byte;
    input reg enable;
    input clk;
    output reg data_out;
    output reg [2:0] index;
);




endmodule
